library verilog;
use verilog.vl_types.all;
entity I2Codec_vlg_vec_tst is
end I2Codec_vlg_vec_tst;
